module Moore_1101_gold(rst, clk, in, out);
input  rst, clk;
input  in;

output reg out;

parameter [2:0] S0=3'd0, S1=3'd1, S2=3'd2, S3=3'd3, S4=3'd4;

reg [2:0] cs, ns;

`protected

    MTI!#As<@w[_*HH**To@T?npnU*#HZn3AE\{37?BZ77i[HnX<$VEVW+~o|)"rJxQ#<*\vHHj},A<
    +sERVp?[G+n~N)&iEYi7JX$Uar="lmBQiQ'~WH$$Y}275jYnlnBo5jT]]>=i2v2Zln^Yo[}~I_gV
    mu^9(qw1C_=>u[2=vn7=5zWRk;kQViUOiGg7aBOZIU~\5;WxV^!,1]v$pp_Ro<3F*~<?-l<}'=Uo
    z\}OI]D=Cu5#YiQD=#*meWAnPKQnuT{jk}#wamsl=T'^3#V_;}a1UAzQRz]~Tnro]PI#Xl{D,U~A
    j]%v3n^5SuqX7]!=7kQiQ;#HQu^B5=j[op{2Bu5&I,a5o?B*ry-s>Qx#TGVT8VO49B1'K;[g
`endprotected

endmodule






 